library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port (
        clk      : in  std_logic;
        endereco : in  unsigned(6 downto 0);   -- 7 bits para 128 endereços
        dado     : out unsigned(18 downto 0)   -- 19 bits de largura
    );
end rom;

architecture a_rom of rom is
    type mem is array (0 to 127) of unsigned(18 downto 0);
    constant conteudo_rom : mem := (
        0  => "0100000000000000001", --LOADAC 1
        1  => "1100000100000000000", --MOVREG R1
        2  => "0000000100000000010", --MOVRAM R1
        3  => "1001000000000000001", --ADDI 1
        4  => "1111000000000100001", --CMPI 33
        5  => "1010000000100000000", --BHI 2
        6  => "0010000000100000000", --JUMP 1
        7  => "0100000000000000100", --LOADAC 4
        8  => "1111000000000100001", --CMPI 33
        9  => "1010000001110000000", --BHI 7
        10 => "1100000100000000000", --MOVREG R1
        11 => "0100000000000000000", --LOADAC 0
        12 => "0000000100000000010", --MOVRAM R1
        13 => "1000000100000000000", --MOVAC R1
        14 => "1001000000000000010", --ADDI 2
        15 => "0010000100000000000", --JUMP 8
        16 => "0100000000000000110", --LOADAC 6
        17 => "1111000000000100001", --CMPI 33
        18 => "1010000001110000000", --BHI 7
        19 => "1100000100000000000", --MOVREG R1
        20 => "0100000000000000000", --LOADAC 0
        21 => "0000000100000000010", --MOVRAM R1
        22 => "1000000100000000000", --MOVAC R1
        23 => "1001000000000000011", --ADDI 3
        24 => "0010001000100000000", --JUMP 17
        25 => "0100000000000001010", --LOADAC 10
        26 => "1111000000000100001", --CMPI 33
        27 => "1010000001110000000", --BHI 7
        28 => "1100000100000000000", --MOVREG R1
        29 => "0100000000000000000", --LOADAC 0
        30 => "0000000100000000010", --MOVRAM R1
        31 => "1000000100000000000", --MOVAC R1
        32 => "1001000000000000101", --ADDI 5
        33 => "0010001101000000000", --JUMP 26
        34 => "0100000000000000001", --LOADAC 1 
        35 => "1111000000000100001", --CMPI 33
        36 => "1010000001110000000", --BHI 7
        37 => "1100000100000000000", --MOVREG R1
        38 => "0000000100000000001", --LOADRAM R1
        39 => "1100001000000000000", --LOADREG R2
        40 => "1000000100000000000", --MOVAC R1
        41 => "1001000000000000001", --ADDI 1
        42 => "0010010001100000000", --JUMP 35
        others => "0000000000000000000"
    );

begin
    process(clk)
    begin
        if rising_edge(clk) then
            dado <= conteudo_rom(to_integer(endereco));
        end if;
    end process;
end architecture;
